.SUBCKT Maxpooling VDD VSS  IN_0[1] IN_0[0] IN_1[1] IN_1[0] IN_2[1] IN_2[0] IN_3[1] IN_3[0] Output[1] Output[0]
XU22 IN_3[1] VDD VSS  n20 INVx8_ASAP7_75t_R
XU23 IN_2[1] VDD VSS  n21 INVx8_ASAP7_75t_R
XU24 IN_1[1] VDD VSS  n22 INVx8_ASAP7_75t_R
XU25 IN_3[1] VDD VSS  n34 INVx8_ASAP7_75t_R
XU26 IN_2[1] VDD VSS  n33 INVx8_ASAP7_75t_R
XU27 IN_1[1] VDD VSS  n42 INVx8_ASAP7_75t_R
XU28 IN_0[1] VDD VSS  n23 INVx8_ASAP7_75t_R
XU29 IN_0[1] VDD VSS  n24 INVx8_ASAP7_75t_R
XU30 IN_0[1] VDD VSS  n41 INVx8_ASAP7_75t_R
XU31 IN_3[1] IN_3[0] VDD VSS  n30 NAND2xp33_ASAP7_75t_R
XU32 n30 IN_1[1] VDD VSS  n32 NAND2xp33_ASAP7_75t_R
XU33 IN_3[1] IN_2[1] VDD VSS  n43 NOR2xp33_ASAP7_75t_R
XU34 n43 IN_0[0] VDD VSS  n29 NAND2xp33_ASAP7_75t_R
XU35 n21 IN_3[0] VDD VSS  n26 NAND2xp33_ASAP7_75t_R
XU36 n20 IN_2[0] VDD VSS  n25 NAND2xp33_ASAP7_75t_R
XU37 n26 n25 VDD VSS  n27 NAND2xp33_ASAP7_75t_R
XU38 n23 n27 VDD VSS  n28 NAND2xp33_ASAP7_75t_R
XU39 n30 n29 n28 VDD VSS  n31 NAND3xp33_ASAP7_75t_R
XU40 n32 n31 VDD VSS  n40 NAND2xp33_ASAP7_75t_R
XU41 n34 n33 n24 VDD VSS  n35 NAND3xp33_ASAP7_75t_R
XU42 n22 n35 VDD VSS  n36 NAND2xp33_ASAP7_75t_R
XU43 IN_1[0] n36 VDD VSS  n39 NAND2xp33_ASAP7_75t_R
XU44 IN_2[1] IN_2[0] VDD VSS  n38 NAND2xp33_ASAP7_75t_R
XU45 IN_0[0] IN_0[1] VDD VSS  n37 NAND2xp33_ASAP7_75t_R
XU46 n40 n39 n38 n37 VDD VSS  Output[0] NAND4xp25_ASAP7_75t_R
XU47 n43 n42 n41 VDD VSS  Output[1] NAND3xp33_ASAP7_75t_R
.ENDS


